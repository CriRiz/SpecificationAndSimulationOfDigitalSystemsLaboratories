
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/21/2025 04:26:16 PM
-- Design Name: 
-- Module Name: Reg - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Reg is
    port(d, d_1, clk, er, rst: IN std_logic;
    q: OUT std_logic);
end Reg;

architecture Behavioral of Reg is

begin
    process(clk)
        begin
            if(rising_edge(clk)) then
                if (rst = '1') then
                    q <= d_1;
                elsif (er = '1') then
                    q <= d;
                end if;
            end if;
    end process;

end Behavioral;
