----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09.10.2025 21:48:14
-- Design Name: 
-- Module Name: Count4to2D - Dataflow
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Count4to2D is
    PORT(d: IN std_logic_vector(3 downto 0);
        q: OUT std_logic_vector(1 downto 0));
end Count4to2D;

architecture Dataflow of Count4to2D is

begin
    q <= "00" when d = "0001" else
    "01" when d = "0010" else
    "10" when d = "0100" else
    "11" when d = "1000" else
    "XX";

end Dataflow;
